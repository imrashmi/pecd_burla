*
.tran 50us 100ms uic
.include rectifier.net

