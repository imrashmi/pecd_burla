*Buck-Boost converter circuit
*
.tran 1us 100ms uic
.include bucboo.net

* Control commands
.control
set color0 = white    	; set background as white
set color1 = black	; set foreground as black
run
plot i(L)
.endc
